library verilog;
use verilog.vl_types.all;
entity atest12 is
end atest12;
