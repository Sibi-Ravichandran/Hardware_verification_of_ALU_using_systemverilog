library verilog;
use verilog.vl_types.all;
entity monitor_sv_unit is
end monitor_sv_unit;
