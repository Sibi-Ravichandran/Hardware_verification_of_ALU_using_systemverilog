library verilog;
use verilog.vl_types.all;
entity adder_test is
end adder_test;
