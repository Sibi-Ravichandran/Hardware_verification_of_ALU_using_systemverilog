library verilog;
use verilog.vl_types.all;
entity A is
end A;
