library verilog;
use verilog.vl_types.all;
entity atest5 is
end atest5;
