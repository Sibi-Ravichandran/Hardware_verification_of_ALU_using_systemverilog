library verilog;
use verilog.vl_types.all;
entity dut_out_c_sv_unit is
end dut_out_c_sv_unit;
