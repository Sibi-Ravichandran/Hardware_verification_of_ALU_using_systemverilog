library verilog;
use verilog.vl_types.all;
entity atest10 is
end atest10;
