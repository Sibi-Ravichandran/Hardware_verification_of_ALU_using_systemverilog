library verilog;
use verilog.vl_types.all;
entity atestreqs is
end atestreqs;
