library verilog;
use verilog.vl_types.all;
entity atest4 is
end atest4;
