library verilog;
use verilog.vl_types.all;
entity driver_sv_unit is
end driver_sv_unit;
