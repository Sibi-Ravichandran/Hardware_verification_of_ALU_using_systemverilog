library verilog;
use verilog.vl_types.all;
entity priority is
    port(
        port1_invalid_op: out    vl_logic;
        port1_invalid_tag: out    vl_logic_vector(0 to 1);
        port2_invalid_op: out    vl_logic;
        port2_invalid_tag: out    vl_logic_vector(0 to 1);
        port3_invalid_op: out    vl_logic;
        port3_invalid_tag: out    vl_logic_vector(0 to 1);
        port4_invalid_op: out    vl_logic;
        port4_invalid_tag: out    vl_logic_vector(0 to 1);
        prio_adder_cmd  : out    vl_logic_vector(0 to 3);
        prio_adder_data1: out    vl_logic_vector(0 to 4);
        prio_adder_data2: out    vl_logic_vector(0 to 4);
        prio_adder_follow_branch: out    vl_logic_vector(0 to 4);
        prio_adder_out_vld: out    vl_logic;
        prio_adder_result: out    vl_logic_vector(0 to 4);
        prio_adder_tag  : out    vl_logic_vector(0 to 3);
        prio_shift_cmd  : out    vl_logic_vector(0 to 3);
        prio_shift_data1: out    vl_logic_vector(0 to 4);
        prio_shift_data2: out    vl_logic_vector(0 to 4);
        prio_shift_data : out    vl_logic_vector(0 to 31);
        prio_shift_follow_branch: out    vl_logic_vector(0 to 4);
        prio_shift_out_vld: out    vl_logic;
        prio_shift_result: out    vl_logic_vector(0 to 4);
        prio_shift_tag  : out    vl_logic_vector(0 to 3);
        scan_out        : out    vl_logic;
        a_clk           : in     vl_logic;
        b_clk           : in     vl_logic;
        c_clk           : in     vl_logic;
        hold1_cmd       : in     vl_logic_vector(0 to 3);
        hold1_data1     : in     vl_logic_vector(0 to 3);
        hold1_data2     : in     vl_logic_vector(0 to 3);
        hold1_data      : in     vl_logic_vector(0 to 31);
        hold1_result    : in     vl_logic_vector(0 to 3);
        hold1_tag       : in     vl_logic_vector(0 to 1);
        hold2_cmd       : in     vl_logic_vector(0 to 3);
        hold2_data1     : in     vl_logic_vector(0 to 3);
        hold2_data2     : in     vl_logic_vector(0 to 3);
        hold2_data      : in     vl_logic_vector(0 to 31);
        hold2_result    : in     vl_logic_vector(0 to 3);
        hold2_tag       : in     vl_logic_vector(0 to 1);
        hold3_cmd       : in     vl_logic_vector(0 to 3);
        hold3_data1     : in     vl_logic_vector(0 to 3);
        hold3_data2     : in     vl_logic_vector(0 to 3);
        hold3_data      : in     vl_logic_vector(0 to 31);
        hold3_result    : in     vl_logic_vector(0 to 3);
        hold3_tag       : in     vl_logic_vector(0 to 1);
        hold4_cmd       : in     vl_logic_vector(0 to 3);
        hold4_data1     : in     vl_logic_vector(0 to 3);
        hold4_data2     : in     vl_logic_vector(0 to 3);
        hold4_data      : in     vl_logic_vector(0 to 31);
        hold4_result    : in     vl_logic_vector(0 to 3);
        hold4_tag       : in     vl_logic_vector(0 to 1);
        reset           : in     vl_logic;
        scan_in         : in     vl_logic
    );
end priority;
