library verilog;
use verilog.vl_types.all;
entity exdbin_mac_test is
end exdbin_mac_test;
