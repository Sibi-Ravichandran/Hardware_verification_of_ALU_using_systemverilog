library verilog;
use verilog.vl_types.all;
entity atest3 is
end atest3;
