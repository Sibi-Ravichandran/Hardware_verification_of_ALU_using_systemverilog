library verilog;
use verilog.vl_types.all;
entity atestsimple is
end atestsimple;
