library verilog;
use verilog.vl_types.all;
entity atest13 is
end atest13;
