library verilog;
use verilog.vl_types.all;
entity atest8 is
end atest8;
