library verilog;
use verilog.vl_types.all;
entity atest1 is
end atest1;
