library verilog;
use verilog.vl_types.all;
entity atest2 is
end atest2;
