library verilog;
use verilog.vl_types.all;
entity atest6and7 is
end atest6and7;
