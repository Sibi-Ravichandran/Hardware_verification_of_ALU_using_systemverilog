library verilog;
use verilog.vl_types.all;
entity atest9 is
end atest9;
