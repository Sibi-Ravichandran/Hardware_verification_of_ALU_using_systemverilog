library verilog;
use verilog.vl_types.all;
entity gen_sv_unit is
end gen_sv_unit;
