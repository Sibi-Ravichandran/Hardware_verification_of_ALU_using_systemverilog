library verilog;
use verilog.vl_types.all;
entity holdreg_test is
end holdreg_test;
