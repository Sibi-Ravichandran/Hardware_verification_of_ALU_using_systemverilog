library verilog;
use verilog.vl_types.all;
entity atest11 is
end atest11;
